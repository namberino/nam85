module top_design(
    input clk
);

    

endmodule
